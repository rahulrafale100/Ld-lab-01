module notgate16(y,x);
output [15:0]y;
input [15:0]x;
notgate notgate_1 [15:0](y,x);
endmodule
